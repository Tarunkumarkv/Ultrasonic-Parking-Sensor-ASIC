module parking_sensor_top (alarm_warning,
    clk,
    echo_pulse,
    reset,
    trigger_pulse);
 output alarm_warning;
 input clk;
 input echo_pulse;
 input reset;
 output trigger_pulse;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire \comp_inst.distance_value[0] ;
 wire \comp_inst.distance_value[10] ;
 wire \comp_inst.distance_value[11] ;
 wire \comp_inst.distance_value[12] ;
 wire \comp_inst.distance_value[13] ;
 wire \comp_inst.distance_value[14] ;
 wire \comp_inst.distance_value[15] ;
 wire \comp_inst.distance_value[1] ;
 wire \comp_inst.distance_value[2] ;
 wire \comp_inst.distance_value[3] ;
 wire \comp_inst.distance_value[4] ;
 wire \comp_inst.distance_value[5] ;
 wire \comp_inst.distance_value[6] ;
 wire \comp_inst.distance_value[7] ;
 wire \comp_inst.distance_value[8] ;
 wire \comp_inst.distance_value[9] ;
 wire \fsm_inst.current_state[0] ;
 wire \fsm_inst.current_state[1] ;
 wire \fsm_inst.current_state[2] ;
 wire \fsm_inst.trigger_done ;
 wire \trig_inst.count[0] ;
 wire \trig_inst.count[1] ;
 wire \trig_inst.count[2] ;
 wire \trig_inst.count[3] ;
 wire \trig_inst.count[4] ;
 wire \trig_inst.count[5] ;
 wire \trig_inst.count[6] ;
 wire \trig_inst.count[7] ;
 wire \trig_inst.count[8] ;
 wire \trig_inst.count[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;

 sky130_fd_sc_hd__inv_2 _115_ (.A(\trig_inst.count[6] ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _116_ (.A(\trig_inst.count[5] ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(net2),
    .Y(_004_));
 sky130_fd_sc_hd__and2_1 _118_ (.A(\comp_inst.distance_value[13] ),
    .B(\comp_inst.distance_value[12] ),
    .X(_114_));
 sky130_fd_sc_hd__and3_1 _119_ (.A(\comp_inst.distance_value[14] ),
    .B(\comp_inst.distance_value[13] ),
    .C(\comp_inst.distance_value[12] ),
    .X(_062_));
 sky130_fd_sc_hd__and4b_2 _120_ (.A_N(net7),
    .B(net11),
    .C(net15),
    .D(net1),
    .X(_063_));
 sky130_fd_sc_hd__and4_1 _121_ (.A(\comp_inst.distance_value[5] ),
    .B(\comp_inst.distance_value[4] ),
    .C(\comp_inst.distance_value[3] ),
    .D(\comp_inst.distance_value[2] ),
    .X(_064_));
 sky130_fd_sc_hd__and4_1 _122_ (.A(\comp_inst.distance_value[7] ),
    .B(\comp_inst.distance_value[6] ),
    .C(\comp_inst.distance_value[1] ),
    .D(\comp_inst.distance_value[0] ),
    .X(_065_));
 sky130_fd_sc_hd__and3_1 _123_ (.A(_063_),
    .B(_064_),
    .C(_065_),
    .X(_066_));
 sky130_fd_sc_hd__and2_1 _124_ (.A(\comp_inst.distance_value[9] ),
    .B(\comp_inst.distance_value[8] ),
    .X(_067_));
 sky130_fd_sc_hd__and4_2 _125_ (.A(_063_),
    .B(_064_),
    .C(_065_),
    .D(_067_),
    .X(_068_));
 sky130_fd_sc_hd__and3_1 _126_ (.A(\comp_inst.distance_value[11] ),
    .B(\comp_inst.distance_value[10] ),
    .C(_068_),
    .X(_069_));
 sky130_fd_sc_hd__and4_1 _127_ (.A(\comp_inst.distance_value[11] ),
    .B(\comp_inst.distance_value[10] ),
    .C(_062_),
    .D(_068_),
    .X(_070_));
 sky130_fd_sc_hd__xor2_1 _128_ (.A(net26),
    .B(_070_),
    .X(_061_));
 sky130_fd_sc_hd__a41o_1 _129_ (.A1(\comp_inst.distance_value[11] ),
    .A2(\comp_inst.distance_value[10] ),
    .A3(_114_),
    .A4(_068_),
    .B1(\comp_inst.distance_value[14] ),
    .X(_071_));
 sky130_fd_sc_hd__and2b_1 _130_ (.A_N(_070_),
    .B(_071_),
    .X(_060_));
 sky130_fd_sc_hd__a41o_1 _131_ (.A1(\comp_inst.distance_value[12] ),
    .A2(\comp_inst.distance_value[11] ),
    .A3(\comp_inst.distance_value[10] ),
    .A4(_068_),
    .B1(\comp_inst.distance_value[13] ),
    .X(_072_));
 sky130_fd_sc_hd__a21boi_1 _132_ (.A1(_114_),
    .A2(_069_),
    .B1_N(_072_),
    .Y(_059_));
 sky130_fd_sc_hd__xor2_1 _133_ (.A(net34),
    .B(_069_),
    .X(_058_));
 sky130_fd_sc_hd__a21oi_1 _134_ (.A1(\comp_inst.distance_value[10] ),
    .A2(_068_),
    .B1(\comp_inst.distance_value[11] ),
    .Y(_073_));
 sky130_fd_sc_hd__nor2_1 _135_ (.A(_069_),
    .B(_073_),
    .Y(_057_));
 sky130_fd_sc_hd__xor2_1 _136_ (.A(net35),
    .B(_068_),
    .X(_056_));
 sky130_fd_sc_hd__a21o_1 _137_ (.A1(\comp_inst.distance_value[8] ),
    .A2(_066_),
    .B1(\comp_inst.distance_value[9] ),
    .X(_074_));
 sky130_fd_sc_hd__and2b_1 _138_ (.A_N(_068_),
    .B(_074_),
    .X(_055_));
 sky130_fd_sc_hd__xor2_1 _139_ (.A(net30),
    .B(_066_),
    .X(_054_));
 sky130_fd_sc_hd__and3_1 _140_ (.A(\comp_inst.distance_value[1] ),
    .B(\comp_inst.distance_value[0] ),
    .C(_063_),
    .X(_075_));
 sky130_fd_sc_hd__and3_1 _141_ (.A(\comp_inst.distance_value[3] ),
    .B(\comp_inst.distance_value[2] ),
    .C(\comp_inst.distance_value[1] ),
    .X(_076_));
 sky130_fd_sc_hd__and3_1 _142_ (.A(\comp_inst.distance_value[0] ),
    .B(_063_),
    .C(_076_),
    .X(_077_));
 sky130_fd_sc_hd__and4_1 _143_ (.A(\comp_inst.distance_value[4] ),
    .B(\comp_inst.distance_value[0] ),
    .C(_063_),
    .D(_076_),
    .X(_078_));
 sky130_fd_sc_hd__and3_1 _144_ (.A(\comp_inst.distance_value[6] ),
    .B(\comp_inst.distance_value[5] ),
    .C(_078_),
    .X(_079_));
 sky130_fd_sc_hd__xor2_1 _145_ (.A(net32),
    .B(_079_),
    .X(_053_));
 sky130_fd_sc_hd__a21oi_1 _146_ (.A1(\comp_inst.distance_value[5] ),
    .A2(_078_),
    .B1(net41),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_1 _147_ (.A(_079_),
    .B(_080_),
    .Y(_052_));
 sky130_fd_sc_hd__xor2_1 _148_ (.A(net39),
    .B(_078_),
    .X(_051_));
 sky130_fd_sc_hd__xor2_1 _149_ (.A(net36),
    .B(_077_),
    .X(_050_));
 sky130_fd_sc_hd__and2_1 _150_ (.A(\comp_inst.distance_value[2] ),
    .B(_075_),
    .X(_081_));
 sky130_fd_sc_hd__o21ba_1 _151_ (.A1(\comp_inst.distance_value[3] ),
    .A2(_081_),
    .B1_N(_077_),
    .X(_049_));
 sky130_fd_sc_hd__nor2_1 _152_ (.A(net40),
    .B(_075_),
    .Y(_082_));
 sky130_fd_sc_hd__nor2_1 _153_ (.A(_081_),
    .B(_082_),
    .Y(_048_));
 sky130_fd_sc_hd__a21oi_1 _154_ (.A1(\comp_inst.distance_value[0] ),
    .A2(_063_),
    .B1(net37),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _155_ (.A(_075_),
    .B(net38),
    .Y(_047_));
 sky130_fd_sc_hd__xor2_1 _156_ (.A(net31),
    .B(_063_),
    .X(_046_));
 sky130_fd_sc_hd__o311ai_2 _157_ (.A1(\trig_inst.count[5] ),
    .A2(\trig_inst.count[4] ),
    .A3(\trig_inst.count[3] ),
    .B1(\trig_inst.count[6] ),
    .C1(\trig_inst.count[7] ),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _158_ (.A(\trig_inst.count[9] ),
    .B(\trig_inst.count[8] ),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_2 _159_ (.A(_084_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__nor3b_4 _160_ (.A(net5),
    .B(net9),
    .C_N(net13),
    .Y(_087_));
 sky130_fd_sc_hd__or3b_1 _161_ (.A(net5),
    .B(net9),
    .C_N(net13),
    .X(_088_));
 sky130_fd_sc_hd__a21o_1 _162_ (.A1(_084_),
    .A2(_085_),
    .B1(_088_),
    .X(_089_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_089_),
    .Y(_000_));
 sky130_fd_sc_hd__and2_1 _164_ (.A(net27),
    .B(_087_),
    .X(_045_));
 sky130_fd_sc_hd__and2_1 _165_ (.A(net28),
    .B(_087_),
    .X(_044_));
 sky130_fd_sc_hd__nand2_1 _166_ (.A(\trig_inst.count[1] ),
    .B(\trig_inst.count[0] ),
    .Y(_090_));
 sky130_fd_sc_hd__and3_1 _167_ (.A(\trig_inst.count[2] ),
    .B(\trig_inst.count[1] ),
    .C(\trig_inst.count[0] ),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__and4_1 _169_ (.A(\trig_inst.count[3] ),
    .B(\trig_inst.count[2] ),
    .C(\trig_inst.count[1] ),
    .D(\trig_inst.count[0] ),
    .X(_093_));
 sky130_fd_sc_hd__inv_2 _170_ (.A(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__nand2_1 _171_ (.A(\trig_inst.count[4] ),
    .B(_093_),
    .Y(_095_));
 sky130_fd_sc_hd__nor4_1 _172_ (.A(_112_),
    .B(_113_),
    .C(_086_),
    .D(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__o21a_1 _173_ (.A1(net33),
    .A2(_096_),
    .B1(_087_),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _174_ (.A(\trig_inst.count[0] ),
    .B(_089_),
    .X(_097_));
 sky130_fd_sc_hd__a41o_1 _175_ (.A1(\trig_inst.count[5] ),
    .A2(\trig_inst.count[4] ),
    .A3(_089_),
    .A4(_093_),
    .B1(\trig_inst.count[6] ),
    .X(_098_));
 sky130_fd_sc_hd__and3b_1 _176_ (.A_N(_096_),
    .B(_098_),
    .C(_087_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _177_ (.A1(\trig_inst.count[4] ),
    .A2(_089_),
    .A3(_093_),
    .B1(\trig_inst.count[5] ),
    .X(_099_));
 sky130_fd_sc_hd__o311a_1 _178_ (.A1(_113_),
    .A2(_000_),
    .A3(_095_),
    .B1(_099_),
    .C1(_087_),
    .X(_041_));
 sky130_fd_sc_hd__a21o_1 _179_ (.A1(_089_),
    .A2(_093_),
    .B1(\trig_inst.count[4] ),
    .X(_100_));
 sky130_fd_sc_hd__o211a_1 _180_ (.A1(_086_),
    .A2(_095_),
    .B1(_100_),
    .C1(_087_),
    .X(_040_));
 sky130_fd_sc_hd__a21o_1 _181_ (.A1(_089_),
    .A2(_091_),
    .B1(\trig_inst.count[3] ),
    .X(_101_));
 sky130_fd_sc_hd__o211a_1 _182_ (.A1(_086_),
    .A2(_094_),
    .B1(_101_),
    .C1(_087_),
    .X(_039_));
 sky130_fd_sc_hd__a31o_1 _183_ (.A1(\trig_inst.count[1] ),
    .A2(\trig_inst.count[0] ),
    .A3(_089_),
    .B1(\trig_inst.count[2] ),
    .X(_102_));
 sky130_fd_sc_hd__o211a_1 _184_ (.A1(_086_),
    .A2(_092_),
    .B1(_102_),
    .C1(_087_),
    .X(_038_));
 sky130_fd_sc_hd__o221a_1 _185_ (.A1(_086_),
    .A2(_090_),
    .B1(_097_),
    .B2(\trig_inst.count[1] ),
    .C1(_087_),
    .X(_037_));
 sky130_fd_sc_hd__nor2_1 _186_ (.A(_086_),
    .B(_088_),
    .Y(_001_));
 sky130_fd_sc_hd__o21ba_1 _187_ (.A1(\trig_inst.count[0] ),
    .A2(_001_),
    .B1_N(_097_),
    .X(_036_));
 sky130_fd_sc_hd__nor2_1 _188_ (.A(\fsm_inst.trigger_done ),
    .B(_088_),
    .Y(_103_));
 sky130_fd_sc_hd__and4bb_1 _189_ (.A_N(net7),
    .B_N(net1),
    .C(net15),
    .D(net11),
    .X(_035_));
 sky130_fd_sc_hd__o21bai_1 _190_ (.A1(net7),
    .A2(net15),
    .B1_N(_063_),
    .Y(_104_));
 sky130_fd_sc_hd__a22o_1 _191_ (.A1(net29),
    .A2(_087_),
    .B1(_104_),
    .B2(net11),
    .X(_034_));
 sky130_fd_sc_hd__or4b_1 _192_ (.A(net7),
    .B(net15),
    .C(net1),
    .D_N(net11),
    .X(_105_));
 sky130_fd_sc_hd__o21a_1 _193_ (.A1(_103_),
    .A2(_104_),
    .B1(_105_),
    .X(_033_));
 sky130_fd_sc_hd__or4_1 _194_ (.A(\comp_inst.distance_value[3] ),
    .B(\comp_inst.distance_value[2] ),
    .C(\comp_inst.distance_value[1] ),
    .D(\comp_inst.distance_value[0] ),
    .X(_106_));
 sky130_fd_sc_hd__or4_1 _195_ (.A(\comp_inst.distance_value[7] ),
    .B(\comp_inst.distance_value[6] ),
    .C(\comp_inst.distance_value[5] ),
    .D(\comp_inst.distance_value[4] ),
    .X(_107_));
 sky130_fd_sc_hd__o311a_1 _196_ (.A1(\comp_inst.distance_value[5] ),
    .A2(\comp_inst.distance_value[4] ),
    .A3(\comp_inst.distance_value[3] ),
    .B1(\comp_inst.distance_value[6] ),
    .C1(\comp_inst.distance_value[7] ),
    .X(_108_));
 sky130_fd_sc_hd__or4_1 _197_ (.A(\comp_inst.distance_value[11] ),
    .B(\comp_inst.distance_value[10] ),
    .C(\comp_inst.distance_value[9] ),
    .D(\comp_inst.distance_value[8] ),
    .X(_109_));
 sky130_fd_sc_hd__or4_1 _198_ (.A(\comp_inst.distance_value[15] ),
    .B(\comp_inst.distance_value[14] ),
    .C(\comp_inst.distance_value[13] ),
    .D(\comp_inst.distance_value[12] ),
    .X(_110_));
 sky130_fd_sc_hd__or3_1 _199_ (.A(_108_),
    .B(_109_),
    .C(_110_),
    .X(_111_));
 sky130_fd_sc_hd__o21ba_1 _200_ (.A1(_106_),
    .A2(_107_),
    .B1_N(_111_),
    .X(net3));
 sky130_fd_sc_hd__o31a_1 _201_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_002_));
 sky130_fd_sc_hd__o31a_1 _202_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_003_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(net2),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(net2),
    .Y(_006_));
 sky130_fd_sc_hd__o31a_1 _205_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_007_));
 sky130_fd_sc_hd__o31a_1 _206_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_008_));
 sky130_fd_sc_hd__o31a_1 _207_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_009_));
 sky130_fd_sc_hd__o31a_1 _208_ (.A1(net7),
    .A2(net11),
    .A3(net15),
    .B1(net19),
    .X(_010_));
 sky130_fd_sc_hd__o31a_1 _209_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_011_));
 sky130_fd_sc_hd__o31a_1 _210_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_012_));
 sky130_fd_sc_hd__o31a_1 _211_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_013_));
 sky130_fd_sc_hd__o31a_1 _212_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_014_));
 sky130_fd_sc_hd__o31a_1 _213_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_015_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_016_));
 sky130_fd_sc_hd__o31a_1 _215_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net19),
    .X(_017_));
 sky130_fd_sc_hd__o31a_1 _216_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__o31a_1 _217_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net19),
    .X(_019_));
 sky130_fd_sc_hd__o31a_1 _218_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net20),
    .X(_020_));
 sky130_fd_sc_hd__o31a_1 _219_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net20),
    .X(_021_));
 sky130_fd_sc_hd__o31a_1 _220_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net20),
    .X(_022_));
 sky130_fd_sc_hd__o31a_1 _221_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net18),
    .X(_023_));
 sky130_fd_sc_hd__o31a_1 _222_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net17),
    .X(_024_));
 sky130_fd_sc_hd__o31a_1 _223_ (.A1(net8),
    .A2(net12),
    .A3(net16),
    .B1(net20),
    .X(_025_));
 sky130_fd_sc_hd__o31a_1 _224_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net18),
    .X(_026_));
 sky130_fd_sc_hd__o31a_1 _225_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_027_));
 sky130_fd_sc_hd__o31a_1 _226_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net17),
    .X(_028_));
 sky130_fd_sc_hd__o31a_1 _227_ (.A1(net5),
    .A2(net9),
    .A3(net13),
    .B1(net17),
    .X(_029_));
 sky130_fd_sc_hd__o31a_1 _228_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net18),
    .X(_030_));
 sky130_fd_sc_hd__o31a_1 _229_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net18),
    .X(_031_));
 sky130_fd_sc_hd__o31a_1 _230_ (.A1(net6),
    .A2(net10),
    .A3(net14),
    .B1(net18),
    .X(_032_));
 sky130_fd_sc_hd__dfrtp_1 _231_ (.CLK(clknet_2_2__leaf_clk),
    .D(_000_),
    .RESET_B(_002_),
    .Q(\fsm_inst.trigger_done ));
 sky130_fd_sc_hd__dfrtp_1 _232_ (.CLK(clknet_2_2__leaf_clk),
    .D(_001_),
    .RESET_B(_003_),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _233_ (.CLK(clknet_2_2__leaf_clk),
    .D(_033_),
    .RESET_B(net19),
    .Q(\fsm_inst.current_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _234_ (.CLK(clknet_2_2__leaf_clk),
    .D(_034_),
    .RESET_B(_005_),
    .Q(\fsm_inst.current_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _235_ (.CLK(clknet_2_2__leaf_clk),
    .D(_035_),
    .RESET_B(_006_),
    .Q(\fsm_inst.current_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _236_ (.CLK(clknet_2_2__leaf_clk),
    .D(_036_),
    .RESET_B(_007_),
    .Q(\trig_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _237_ (.CLK(clknet_2_2__leaf_clk),
    .D(_037_),
    .RESET_B(_008_),
    .Q(\trig_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _238_ (.CLK(clknet_2_2__leaf_clk),
    .D(_038_),
    .RESET_B(_009_),
    .Q(\trig_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _239_ (.CLK(clknet_2_2__leaf_clk),
    .D(_039_),
    .RESET_B(_010_),
    .Q(\trig_inst.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _240_ (.CLK(clknet_2_0__leaf_clk),
    .D(_040_),
    .RESET_B(_011_),
    .Q(\trig_inst.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _241_ (.CLK(clknet_2_0__leaf_clk),
    .D(_041_),
    .RESET_B(_012_),
    .Q(\trig_inst.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _242_ (.CLK(clknet_2_0__leaf_clk),
    .D(_042_),
    .RESET_B(_013_),
    .Q(\trig_inst.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _243_ (.CLK(clknet_2_0__leaf_clk),
    .D(_043_),
    .RESET_B(_014_),
    .Q(\trig_inst.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _244_ (.CLK(clknet_2_0__leaf_clk),
    .D(_044_),
    .RESET_B(_015_),
    .Q(\trig_inst.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _245_ (.CLK(clknet_2_0__leaf_clk),
    .D(_045_),
    .RESET_B(_016_),
    .Q(\trig_inst.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _246_ (.CLK(clknet_2_3__leaf_clk),
    .D(_046_),
    .RESET_B(_017_),
    .Q(\comp_inst.distance_value[0] ));
 sky130_fd_sc_hd__dfrtp_1 _247_ (.CLK(clknet_2_3__leaf_clk),
    .D(_047_),
    .RESET_B(net24),
    .Q(\comp_inst.distance_value[1] ));
 sky130_fd_sc_hd__dfrtp_1 _248_ (.CLK(clknet_2_3__leaf_clk),
    .D(_048_),
    .RESET_B(_019_),
    .Q(\comp_inst.distance_value[2] ));
 sky130_fd_sc_hd__dfrtp_1 _249_ (.CLK(clknet_2_3__leaf_clk),
    .D(_049_),
    .RESET_B(_020_),
    .Q(\comp_inst.distance_value[3] ));
 sky130_fd_sc_hd__dfrtp_1 _250_ (.CLK(clknet_2_3__leaf_clk),
    .D(_050_),
    .RESET_B(_021_),
    .Q(\comp_inst.distance_value[4] ));
 sky130_fd_sc_hd__dfrtp_1 _251_ (.CLK(clknet_2_3__leaf_clk),
    .D(_051_),
    .RESET_B(net22),
    .Q(\comp_inst.distance_value[5] ));
 sky130_fd_sc_hd__dfrtp_1 _252_ (.CLK(clknet_2_1__leaf_clk),
    .D(_052_),
    .RESET_B(_023_),
    .Q(\comp_inst.distance_value[6] ));
 sky130_fd_sc_hd__dfrtp_1 _253_ (.CLK(clknet_2_1__leaf_clk),
    .D(_053_),
    .RESET_B(_024_),
    .Q(\comp_inst.distance_value[7] ));
 sky130_fd_sc_hd__dfrtp_1 _254_ (.CLK(clknet_2_3__leaf_clk),
    .D(_054_),
    .RESET_B(_025_),
    .Q(\comp_inst.distance_value[8] ));
 sky130_fd_sc_hd__dfrtp_1 _255_ (.CLK(clknet_2_1__leaf_clk),
    .D(_055_),
    .RESET_B(_026_),
    .Q(\comp_inst.distance_value[9] ));
 sky130_fd_sc_hd__dfrtp_2 _256_ (.CLK(clknet_2_1__leaf_clk),
    .D(_056_),
    .RESET_B(_027_),
    .Q(\comp_inst.distance_value[10] ));
 sky130_fd_sc_hd__dfrtp_1 _257_ (.CLK(clknet_2_1__leaf_clk),
    .D(_057_),
    .RESET_B(_028_),
    .Q(\comp_inst.distance_value[11] ));
 sky130_fd_sc_hd__dfrtp_1 _258_ (.CLK(clknet_2_1__leaf_clk),
    .D(_058_),
    .RESET_B(_029_),
    .Q(\comp_inst.distance_value[12] ));
 sky130_fd_sc_hd__dfrtp_1 _259_ (.CLK(clknet_2_1__leaf_clk),
    .D(_059_),
    .RESET_B(_030_),
    .Q(\comp_inst.distance_value[13] ));
 sky130_fd_sc_hd__dfrtp_1 _260_ (.CLK(clknet_2_1__leaf_clk),
    .D(_060_),
    .RESET_B(_031_),
    .Q(\comp_inst.distance_value[14] ));
 sky130_fd_sc_hd__dfrtp_1 _261_ (.CLK(clknet_2_1__leaf_clk),
    .D(_061_),
    .RESET_B(_032_),
    .Q(\comp_inst.distance_value[15] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(echo_pulse),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(reset),
    .X(net2));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(alarm_warning));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(trigger_pulse));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net25),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 fanout6 (.A(net25),
    .X(net6));
 sky130_fd_sc_hd__buf_2 fanout7 (.A(net25),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 fanout8 (.A(net25),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net23),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 fanout10 (.A(net23),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net23),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net23),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net21),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net21),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net21),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net21),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net20),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout18 (.A(net20),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(_004_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\fsm_inst.current_state[0] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_022_),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\fsm_inst.current_state[1] ),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_018_),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\fsm_inst.current_state[2] ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\comp_inst.distance_value[15] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\trig_inst.count[9] ),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\trig_inst.count[8] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fsm_inst.trigger_done ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\comp_inst.distance_value[8] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\comp_inst.distance_value[0] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\comp_inst.distance_value[7] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\trig_inst.count[7] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\comp_inst.distance_value[12] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\comp_inst.distance_value[10] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\comp_inst.distance_value[4] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\comp_inst.distance_value[1] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_083_),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\comp_inst.distance_value[5] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\comp_inst.distance_value[2] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\comp_inst.distance_value[6] ),
    .X(net41));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_137 ();
endmodule
